/* 
 * Do not change Module name 
*/
module main;
  initial 
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule